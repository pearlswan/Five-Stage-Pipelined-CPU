module DE1_SoC(clk, rst, regw, read1, read2, wdata, data1, data2);
	input clk, rst, regw;
	input [4:0] read1, read2;
	input [63:0] wdata;
	output [63:0] data1, data2;
	
	
endmodule
